b0VIM 7.4      m�e[�$<��  fengmao                                 amax                                    ~fengmao/Adapt_seg/result_IN.txt                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   3210    #"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 tp           f                     ��������g       g                     e       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ad      �     f       �  �  �  v  S  0    �  �  �  �  ^  ;    �  �  �  �  i  F  #     �  �  �  p  L  (    �  �  �  t  P  ,    �
  �
  �
  x
  T
  0
  
  �	  �	  �	  |	  X	  4	  	  �  �  �  �  \  8    �  �  �  �  `  <    �  �  �  �  d  @    �  �  �  �  h  D     �  �  �  �  q  N  +    �  �  �  |  Y  6    �  �  �  �  d  @    �  �  �                                  i_iter:11500,        miou:32.22000  i_iter:11000,        miou:32.55000  i_iter:10500,        miou:32.15000  i_iter:10000,        miou:31.61000  i_iter:9500,        miou:32.10000  i_iter:9000,        miou:32.42000  i_iter:8500,        miou:32.21000  i_iter:8000,        miou:31.92000  i_iter:7500,        miou:31.93000  i_iter:7000,        miou:32.35000  i_iter:6500,        miou:31.51000  i_iter:6000,        miou:31.82000  i_iter:5500,        miou:32.10000  i_iter:5000,        miou:32.02000  i_iter:4500,        miou:30.82000  i_iter:4000,        miou:30.99000  i_iter:3500,        miou:31.15000  i_iter:3000,        miou:30.89000  i_iter:2500,        miou:31.02000  i_iter:2000,        miou:30.75000  i_iter:1500,        miou:30.74000  i_iter:1000,        miou:28.20000  i_iter:500,        miou:26.95000  i_iter:38000,        miou:33.39000  i_iter:37500,        miou:33.07000  i_iter:37000,        miou:33.73000  i_iter:36500,        miou:34.21000  i_iter:36000,        miou:33.80000  i_iter:35500,        miou:33.67000  i_iter:35000,        miou:33.59000  i_iter:34500,        miou:32.82000  i_iter:34000,        miou:32.87000  i_iter:33500,        miou:33.75000  i_iter:33000,        miou:33.32000  i_iter:32500,        miou:33.00000  i_iter:32000,        miou:33.24000  i_iter:31500,        miou:33.10000  i_iter:31000,        miou:33.17000  i_iter:30500,        miou:32.26000  i_iter:30000,        miou:32.70000  i_iter:29500,        miou:32.97000  i_iter:29000,        miou:33.51000  i_iter:28500,        miou:32.74000  i_iter:28000,        miou:32.75000  i_iter:27500,        miou:33.43000  i_iter:27000,        miou:33.01000  i_iter:26500,        miou:32.52000  i_iter:26000,        miou:32.64000  i_iter:25500,        miou:32.67000  i_iter:25000,        miou:32.42000  i_iter:24500,        miou:32.97000  i_iter:24000,        miou:33.02000  i_iter:23500,        miou:32.06000  i_iter:23000,        miou:32.72000  i_iter:22500,        miou:32.75000  i_iter:22000,        miou:33.03000  i_iter:21500,        miou:32.61000  i_iter:21000,        miou:32.76000  i_iter:20500,        miou:32.85000  i_iter:20000,        miou:31.24000  i_iter:19500,        miou:32.15000  i_iter:19000,        miou:32.85000  i_iter:18500,        miou:31.93000  i_iter:18000,        miou:31.78000  i_iter:17500,        miou:32.25000  i_iter:17000,        miou:31.17000  i_iter:16500,        miou:31.44000  i_iter:16000,        miou:32.61000  i_iter:15500,        miou:32.48000  i_iter:15000,        miou:32.60000  i_iter:14500,        miou:32.24000  i_iter:14000,        miou:32.60000  i_iter:13500,        miou:32.84000  i_iter:13000,        miou:32.13000  i_iter:12500,        miou:32.71000  i_iter:12000,        miou:32.88000  i_iter:11500,        miou:32.46000  i_iter:11000,        miou:31.92000  i_iter:10500,        miou:33.09000  i_iter:10000,        miou:32.22000  i_iter:9500,        miou:32.26000  i_iter:9000,        miou:31.97000  i_iter:8500,        miou:32.67000  i_iter:8000,        miou:31.62000  i_iter:7500,        miou:32.20000  i_iter:7000,        miou:31.74000  i_iter:6500,        miou:33.17000  i_iter:6000,        miou:32.25000  i_iter:5500,        miou:32.09000  i_iter:5000,        miou:32.27000  i_iter:4500,        miou:31.75000  i_iter:4000,        miou:31.32000  i_iter:3500,        miou:31.89000  i_iter:3000,        miou:30.65000  i_iter:2500,        miou:30.53000  i_iter:2000,        miou:30.73000  i_iter:1500,        miou:29.59000  i_iter:1000,        miou:27.62000  i_iter:500,        miou:26.93000  i_iter:1500,        miou:29.14000  i_iter:1000,        miou:27.98000  i_iter:500,        miou:27.61000  ad  %   �     e       �  �  �  t  Q  .    �  �  �  }  Y  5    �  �  �  �  ]  9    �  �  �  �  a  =    �  �  �  �  e  A    �
  �
  �
  �
  i
  E
  !
  �	  �	  �	  �	  m	  I	  %	  	  �  �  �  q  M  )    �  �  �  u  Q  -  	  �  �  �  y  U  1    �  �  �  }  Y  5    �  �  �  �  ]  9    �  �  �  �  a  =    �  �  �  �  e  A    �  �  �                                       i_iter:55500,        miou:35.21000  i_iter:55000,        miou:35.02000  i_iter:54500,        miou:36.09000  i_iter:54000,        miou:36.52000  i_iter:53500,        miou:35.21000  i_iter:53000,        miou:33.24000  i_iter:52500,        miou:34.52000  i_iter:52000,        miou:37.20000  i_iter:51500,        miou:33.29000  i_iter:51000,        miou:34.85000  i_iter:50500,        miou:33.72000  i_iter:50000,        miou:34.31000  i_iter:49500,        miou:32.70000  i_iter:49000,        miou:33.76000  i_iter:48500,        miou:33.66000  i_iter:48000,        miou:32.36000  i_iter:47500,        miou:30.65000  i_iter:47000,        miou:29.65000  i_iter:46500,        miou:32.04000  i_iter:46000,        miou:32.23000  i_iter:45500,        miou:32.73000  i_iter:45000,        miou:32.00000  i_iter:44500,        miou:32.18000  i_iter:44000,        miou:34.98000  i_iter:43500,        miou:31.87000  i_iter:43000,        miou:32.81000  i_iter:42500,        miou:33.39000  i_iter:42000,        miou:34.81000  i_iter:41500,        miou:34.46000  i_iter:41000,        miou:35.64000  i_iter:40500,        miou:34.58000  i_iter:40000,        miou:33.58000  i_iter:39500,        miou:34.83000  i_iter:39000,        miou:33.25000  i_iter:38500,        miou:36.41000  i_iter:38000,        miou:32.18000  i_iter:37500,        miou:30.80000  i_iter:37000,        miou:34.90000  i_iter:36500,        miou:34.94000  i_iter:36000,        miou:32.23000  i_iter:35500,        miou:31.86000  i_iter:35000,        miou:31.57000  i_iter:34500,        miou:34.04000  i_iter:34000,        miou:34.08000  i_iter:33500,        miou:37.50000  i_iter:33000,        miou:32.99000  i_iter:32500,        miou:32.42000  i_iter:32000,        miou:33.04000  i_iter:31500,        miou:36.62000  i_iter:31000,        miou:30.82000  i_iter:30500,        miou:34.17000  i_iter:30000,        miou:32.86000  i_iter:29500,        miou:30.58000  i_iter:29000,        miou:31.54000  i_iter:28500,        miou:34.19000  i_iter:28000,        miou:32.25000  i_iter:27500,        miou:32.09000  i_iter:27000,        miou:33.24000  i_iter:26500,        miou:31.70000  i_iter:26000,        miou:35.26000  i_iter:25500,        miou:29.34000  i_iter:25000,        miou:31.93000  i_iter:24500,        miou:32.36000  i_iter:24000,        miou:31.55000  i_iter:23500,        miou:31.17000  i_iter:23000,        miou:31.36000  i_iter:22500,        miou:33.13000  i_iter:22000,        miou:28.63000  i_iter:21500,        miou:31.37000  i_iter:21000,        miou:31.35000  i_iter:20500,        miou:31.02000  i_iter:20000,        miou:31.53000  i_iter:19500,        miou:30.83000  i_iter:19000,        miou:31.17000  i_iter:18500,        miou:34.12000  i_iter:18000,        miou:32.48000  i_iter:17500,        miou:31.40000  i_iter:17000,        miou:31.65000  i_iter:16500,        miou:31.00000  i_iter:16000,        miou:30.77000  i_iter:15500,        miou:31.79000  i_iter:15000,        miou:34.27000  i_iter:14500,        miou:31.17000  i_iter:14000,        miou:30.12000  i_iter:13500,        miou:30.68000  i_iter:13000,        miou:28.75000  i_iter:12500,        miou:31.18000  i_iter:12000,        miou:30.87000  i_iter:11500,        miou:28.22000  i_iter:11000,        miou:31.35000  i_iter:10500,        miou:29.49000  i_iter:10000,        miou:28.47000  i_iter:9500,        miou:29.76000  i_iter:9000,        miou:29.38000  i_iter:8500,        miou:29.26000  i_iter:8000,        miou:27.09000  i_iter:7500,        miou:30.81000  i_iter:7000,        miou:28.49000  i_iter:6500,        miou:30.28000  i_iter:6000,        miou:28.92000  i_iter:5500,        miou:29.17000  