b0VIM 7.4      �f[�$<JO  fengmao                                 amax                                    ~fengmao/Adapt_seg/result_lse_drop.txt                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             3210    #"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 tp           g                     ��������f       h                            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ad     �     g       �  �  �  u  R  /    �  �  �  �  ]  :    �  �  �  �  h  D     �  �  �  �  l  H  $     �  �  �  p  L  (    �
  �
  �
  t
  P
  ,
  
  �	  �	  �	  x	  T	  0	  	  �  �  �  |  X  4    �  �  �  �  \  :    �  �  �  �  h  E  "  �  �  �  �  s  P  -  
  �  �  �  ~  [  9    �  �  �  �  h  E  "  �  �  �  �  u  R  /    �  �  �                i_iter:3000,        miou:32.79000  i_iter:2500,        miou:36.58000  i_iter:2000,        miou:36.85000  i_iter:1500,        miou:33.36000  i_iter:1000,        miou:25.71000  i_iter:500,        miou:27.56000  i_iter:500,        miou:24.26000  i_iter:5000,        miou:34.08000  i_iter:4500,        miou:36.68000  i_iter:4000,        miou:34.45000  i_iter:3500,        miou:36.68000  i_iter:3000,        miou:36.25000  i_iter:2500,        miou:34.79000  i_iter:2000,        miou:34.85000  i_iter:1500,        miou:32.65000  i_iter:1000,        miou:29.44000  i_iter:500,        miou:26.21000  i_iter:1000,        miou:28.43000  i_iter:500,        miou:25.98000  i_iter:1000,        miou:22.83000  i_iter:500,        miou:20.85000  i_iter:10000,        miou:36.15000  i_iter:9500,        miou:37.38000  i_iter:9000,        miou:40.65000  i_iter:8500,        miou:36.46000  i_iter:8000,        miou:41.99000  i_iter:7500,        miou:41.17000  i_iter:7000,        miou:37.76000  i_iter:6500,        miou:40.99000  i_iter:6000,        miou:40.00000  i_iter:5500,        miou:42.67000  i_iter:5000,        miou:40.13000  i_iter:4500,        miou:42.13000  i_iter:4000,        miou:40.01000  i_iter:3500,        miou:36.96000  i_iter:3000,        miou:37.78000  i_iter:2500,        miou:38.12000  i_iter:2000,        miou:38.25000  i_iter:1500,        miou:38.53000  i_iter:1000,        miou:36.90000  i_iter:500,        miou:37.10000  i_iter:31000,        miou:44.79000  i_iter:30500,        miou:44.75000  i_iter:30000,        miou:43.65000  i_iter:29500,        miou:42.61000  i_iter:29000,        miou:44.61000  i_iter:28500,        miou:44.49000  i_iter:28000,        miou:44.80000  i_iter:27500,        miou:44.25000  i_iter:27000,        miou:44.37000  i_iter:26500,        miou:44.98000  i_iter:26000,        miou:44.22000  i_iter:25500,        miou:44.96000  i_iter:25000,        miou:43.32000  i_iter:24500,        miou:44.23000  i_iter:24000,        miou:44.75000  i_iter:23500,        miou:44.88000  i_iter:23000,        miou:43.60000  i_iter:22500,        miou:43.77000  i_iter:22000,        miou:43.56000  i_iter:21500,        miou:44.18000  i_iter:21000,        miou:44.94000  i_iter:20500,        miou:42.59000  i_iter:20000,        miou:41.68000  i_iter:19500,        miou:44.73000  i_iter:19000,        miou:43.98000  i_iter:18500,        miou:43.60000  i_iter:18000,        miou:44.98000  i_iter:17500,        miou:45.14000  i_iter:17000,        miou:44.21000  i_iter:16500,        miou:43.45000  i_iter:16000,        miou:43.35000  i_iter:15500,        miou:43.49000  i_iter:15000,        miou:42.35000  i_iter:14500,        miou:43.53000  i_iter:14000,        miou:43.07000  i_iter:13500,        miou:42.70000  i_iter:13000,        miou:42.29000  i_iter:12500,        miou:43.89000  i_iter:12000,        miou:41.36000  i_iter:11500,        miou:42.85000  i_iter:11000,        miou:44.27000  i_iter:10500,        miou:43.29000  i_iter:10000,        miou:42.04000  i_iter:9500,        miou:42.30000  i_iter:9000,        miou:42.60000  i_iter:8500,        miou:42.10000  i_iter:8000,        miou:41.57000  i_iter:7500,        miou:41.42000  i_iter:7000,        miou:42.85000  i_iter:6500,        miou:40.05000  i_iter:6000,        miou:41.63000  i_iter:5500,        miou:40.19000  i_iter:5000,        miou:39.68000  i_iter:4500,        miou:39.78000  i_iter:4000,        miou:39.01000  i_iter:3500,        miou:39.02000  i_iter:3000,        miou:38.30000  i_iter:2500,        miou:35.78000  i_iter:2000,        miou:37.00000  i_iter:1500,        miou:32.82000  i_iter:1000,        miou:32.93000  i_iter:500,        miou:29.85000  ad  t  �            �  �  �  p  L  (    �  �  �  t  P  ,    �  �  �  x  T  0    �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      i_iter:65500,        miou:46.20000  i_iter:65000,        miou:47.13000  i_iter:64500,        miou:46.06000  i_iter:63500,        miou:44.97000  i_iter:63000,        miou:41.87000  i_iter:62500,        miou:44.19000  i_iter:62000,        miou:45.22000  i_iter:61500,        miou:44.15000  i_iter:61000,        miou:45.53000  i_iter:60500,        miou:45.00000  i_iter:60000,        miou:42.69000  i_iter:59500,        miou:43.83000  i_iter:59000,        miou:41.44000  i_iter:58500,        miou:41.07000  i_iter:58000,        miou:44.46000  i_iter:57500,        miou:43.72000  i_iter:57000,        miou:41.01000  i_iter:56500,        miou:43.75000  i_iter:56000,        miou:43.15000  i_iter:55500,        miou:42.76000  i_iter:55000,        miou:42.98000  i_iter:54500,        miou:43.76000  